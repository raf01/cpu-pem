module acumulador();

endmodule