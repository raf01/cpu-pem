module registrador(operando);
input [7:0]operando;

endmodule

